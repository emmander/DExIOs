module andGate(
	input wire a,b,
	output wire q
	);
	assign q = a & b;
	endmodule